`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05.01.2024 14:44:43
// Design Name: 
// Module Name: FULL_SUBTRACTOR
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module full_subtractor(a, b, c, D, Bout);
input a, b, c;
output D, Bout;
assign D = a ^ b ^ c ;
assign Bout = ~a & (b^c) | b & c;
endmodule
